netcdf glider_trajectory_v.0.0 {
dimensions:
	trajectory = 1 ;
    time_avg = 1 ;
	time = 1076 ;
variables:
	int trajectory(trajectory) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:long_name = "Unique identifier for each trajectory feature instance" ;
	double time(time) ;
		time:axis = "T" ;
		time:calendar = "gregorian" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;
	double time_avg(time_avg) ;
		time_avg:axis = "T" ;
		time_avg:calendar = "gregorian" ;
		time_avg:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time_avg:standard_name = "time" ;
		time_avg:long_name = "Time corresponding to midpoint of segment" ;
		time_avg:observation_type = "measured" ;
	int segment_id(time) ;
		segment_id:_FillValue = -2147483647 ;
		segment_id:comment = "Sequential segment number for the trajectory.  A segment is defined the collection of profiles contained in the trajectory" ;
		segment_id:long_name = "Segment ID" ;
		segment_id:valid_min = 1 ;
		segment_id:valid_max = 999 ;
		segment_id:observation_type = "calculated" ;
		segment_id:ancillary_variables = "slocum profile_id trajectory" ;
		segment_id:platform = "slocum" ;
	int profile_id(time) ;
		profile_id:_FillValue = -2147483647 ;
		profile_id:comment = "Sequential profile number contained in the trajectory.  A profile is defined a single dive or climb" ;
		profile_id:long_name = "Profile ID" ;
		profile_id:valid_min = 1 ;
		profile_id:valid_max = 999 ;
		profile_id:observation_type = "calculated" ;
		profile_id:ancillary_variables = "slocum segment_id trajectory" ;
		profile_id:platform = "slocum" ;
	double depth(time) ;
		depth:_FillValue = 9.96920996838687e+36 ;
		depth:axis = "Z" ;
		depth:units = "meters" ;
		depth:standard_name = "depth" ;
		depth:valid_min = 0. ;
		depth:valid_max = 2000. ;
		depth:long_name = "Depth" ;
		depth:reference_datum = "sea-surface" ;
		depth:vertical_positive = "down" ;
		depth:observation_type = "calculated" ;
		depth:ancillary_variables = "depth_qc instrument_ctd" ;
		depth:platform = "slocum" ;
		depth:instrument = "instrument_ctd" ;
	byte depth_qc(time) ;
		depth_qc:_FillValue = -127b ;
		depth_qc:long_name = "depth Quality" ;
		depth_qc:standard_name = "depth status_flag" ;
		depth_qc:flag_meanings = "" ;
		depth_qc:valid_range = 0., 128. ;
		depth_qc:flag_values = "" ;
		depth_qc:ancillary_variables = "depth instrument_ctd" ;
	double lat(time) ;
		lat:_FillValue = 9.96920996838687e+36 ;
		lat:axis = "Y" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
		lat:long_name = "Latitude" ;
		lat:observation_type = "measured" ;
		lat:ancillary_variables = "lat_qc" ;
		lat:platform = "slocum" ;
	byte lat_qc(time) ;
		lat_qc:_FillValue = -127b ;
		lat_qc:long_name = "lat Quality" ;
		lat_qc:standard_name = "lat status_flag" ;
		lat_qc:flag_meanings = "" ;
		lat_qc:valid_range = 0., 128. ;
		lat_qc:flag_values = "" ;
		lat_qc:ancillary_variables = "lat" ;
	double lon(time) ;
		lon:_FillValue = 9.96920996838687e+36 ;
		lon:axis = "X" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:long_name = "Longitude" ;
		lon:observation_type = "measured" ;
		lon:ancillary_variables = "lon" ;
		lon:platform = "slocum" ;
	byte lon_qc(time) ;
		lon_qc:_FillValue = -127b ;
		lon_qc:long_name = "lon Quality" ;
		lon_qc:standard_name = "lon status_flag" ;
		lon_qc:flag_meanings = "" ;
		lon_qc:valid_range = 0., 128. ;
		lon_qc:flag_values = "" ;
		lon_qc:ancillary_variables = "lon" ;
	double pressure(time) ;
		pressure:_FillValue = 9.96920996838687e+36 ;
		pressure:axis = "Z" ;
		pressure:units = "dbar" ;
		pressure:standard_name = "pressure" ;
		pressure:valid_min = 0. ;
		pressure:valid_max = 2000. ;
		pressure:long_name = "Pressure" ;
		pressure:reference_datum = "sea-surface" ;
		pressure:vertical_positive = "down" ;
		pressure:observation_type = "measured" ;
		pressure:ancillary_variables = "pressure_qc instrument_ctd" ;
		pressure:platform = "slocum" ;
		pressure:instrument = "instrument_ctd" ;
	byte pressure_qc(time) ;
		pressure_qc:_FillValue = -127b ;
		pressure_qc:long_name = "pressure Quality" ;
		pressure_qc:standard_name = "pressure status_flag" ;
		pressure_qc:flag_meanings = "" ;
		pressure_qc:valid_range = 0., 128. ;
		pressure_qc:flag_values = "" ;
		pressure_qc:ancillary_variables = "pressure instrument_ctd" ;
	double conductivity(time) ;
		conductivity:_FillValue = 9.96920996838687e+36 ;
		conductivity:units = "S m-1" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:valid_min = 0. ;
		conductivity:valid_max = 10. ;
		conductivity:long_name = "Sea Water Conductivity" ;
		conductivity:observation_type = "measured" ;
		conductivity:coordinates = "lon lat depth time" ;
		conductivity:ancillary_variables = "conductivity instrument_ctd" ;
		conductivity:platform = "slocum" ;
		conductivity:instrument = "instrument_ctd" ;
	byte conductivity_qc(time) ;
		conductivity_qc:_FillValue = -127b ;
		conductivity_qc:long_name = "conductivity Quality" ;
		conductivity_qc:standard_name = "conductivity status_flag" ;
		conductivity_qc:flag_meanings = "" ;
		conductivity_qc:valid_range = 0., 128. ;
		conductivity_qc:flag_values = "" ;
	double density(time) ;
		density:_FillValue = 9.96920996838687e+36 ;
		density:units = "kg m-3" ;
		density:standard_name = "sea_water_density" ;
		density:valid_min = 1015. ;
		density:valid_max = 1040. ;
		density:long_name = "Sea Water Density" ;
		density:observation_type = "calculated" ;
		density:coordinates = "lon lat depth time" ;
		density:ancillary_variables = "density_qc instrument_ctd" ;
		density:platform = "slocum" ;
		density:instrument = "instrument_ctd" ;
	byte density_qc(time) ;
		density_qc:_FillValue = -127b ;
		density_qc:long_name = "density Quality" ;
		density_qc:standard_name = "density status_flag" ;
		density_qc:flag_meanings = "" ;
		density_qc:valid_range = 0., 128. ;
		density_qc:flag_values = "" ;
		density_qc:ancillary_variables = "density instrument_ctd" ;
	double salinity(time) ;
		salinity:_FillValue = 9.96920996838687e+36 ;
		salinity:units = "1e-3" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:valid_min = 0. ;
		salinity:valid_max = 40. ;
		salinity:long_name = "Sea Water Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:coordinates = "lon lat depth time" ;
		salinity:ancillary_variables = "salinity_qc instrument_ctd" ;
		salinity:platform = "slocum" ;
		salinity:instrument = "instrument_ctd" ;
	byte salinity_qc(time) ;
		salinity_qc:_FillValue = -127b ;
		salinity_qc:long_name = "salinity Quality" ;
		salinity_qc:standard_name = "salinity status_flag" ;
		salinity_qc:flag_meanings = "" ;
		salinity_qc:valid_range = 0., 128. ;
		salinity_qc:flag_values = "" ;
		salinity_qc:ancillary_variables = "salinity instrument_ctd" ;
	double temperature(time) ;
		temperature:_FillValue = 9.96920996838687e+36 ;
		temperature:units = "Celsius" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:valid_min = -5. ;
		temperature:valid_max = 40. ;
		temperature:long_name = "Sea Water Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:coordinates = "lon lat depth time" ;
		temperature:ancillary_variables = "temperature_qc instrument_ctd" ;
		temperature:platform = "slocum" ;
		temperature:instrument = "instrument_ctd" ;
	byte temperature_qc(time) ;
		temperature_qc:_FillValue = -127b ;
		temperature_qc:long_name = "temperature Quality" ;
		temperature_qc:standard_name = "temperature status_flag" ;
		temperature_qc:flag_meanings = "" ;
		temperature_qc:valid_range = 0., 128. ;
		temperature_qc:flag_values = "" ;
		temperature_qc:ancillary_variables = "temperature instrument_ctd" ;
	double u(time_avg) ;
		u:_FillValue = 9.96920996838687e+36 ;
		u:units = "m s-1" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:valid_min = 0. ;
		u:valid_max = 3. ;
		u:long_name = "Eastward Sea Water Velocity" ;
		u:observation_type = "calculated" ;
		u:coordinates = "time_avg" ;
	byte u_qc(time_avg) ;
		u_qc:_FillValue = -127b ;
		u_qc:long_name = "u Quality" ;
		u_qc:flag_meanings = "" ;
		u_qc:valid_range = 0., 128. ;
		u_qc:flag_values = "" ;
		u_qc:ancillary_variables = "u" ;
	double v(time_avg) ;
		v:_FillValue = 9.96920996838687e+36 ;
		v:units = "m s-1" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:valid_min = 0. ;
		v:valid_max = 3. ;
		v:long_name = "Northward Sea Water Velocity" ;
		v:observation_type = "calculated" ;
		v:coordinates = "time_avg" ;
	byte v_qc(time_avg) ;
		v_qc:_FillValue = -127b ;
		v_qc:long_name = "v Quality" ;
		v_qc:flag_meanings = "" ;
		v_qc:valid_range = 0., 128. ;
		v_qc:flag_values = "" ;
		v_qc:ancillary_variables = "v" ;
	int slocum ;
		slocum:wmo_id = "ru29" ;
		slocum:comment = "Slocum Glider ru29" ;
		slocum:id = "ru29" ;
		slocum:long_name = "Slocum Glider ru29" ;
	int instrument_ctd ;
		instrument_ctd:comment = "Unpumped CTD with a nominal sampling rate of 1Hz." ;
		instrument_ctd:serial_number = -1 ;
		instrument_ctd:long_name = "Seabird SBD 41CP Conductivity, Temperature, Depth Sensor." ;
		instrument_ctd:ancillary_variables = "slocum temperature temperature_qc salinity salinity_qc pressure pressure_qc depth depth_qc conductivity conductivity_qc" ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:acknowledgment = "" ;
        :cdl_template_version = "IOOS_Glider_NetCDF_Trajectory_Template_v0.0" ;
		:cdm_data_type = "Trajectory" ;
		:comment = "" ;
		:contributor_name = "Scott Glenn, Oscar Schofield, John Kerfoot" ;
		:contributor_role = "Principal Investigator, Principal Investigator, Data Manager" ;
		:creator_email = "kerfoot@marine.rutgers.edu" ;
		:creator_name = "John Kerfoot" ;
		:creator_url = "http://marine.rutgers.edu/cool/auvs" ;
		:date_created = "2013-05-08 14:45 UTC" ;
		:date_issued = "2013-05-08 14:45 UTC" ;
		:date_modified = "2013-05-08 14:45 UTC" ;
		:featureType = "trajectory" ;
		:geospatial_lat_max = -15.88833 ;
		:geospatial_lat_min = -15.9445416666667 ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 1.49547333333333 ;
		:geospatial_lon_min = 1.394655 ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_max = 987.26 ;
		:geospatial_vertical_min = 0. ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_units = "meters" ;
		:history = "Created with the Matlab 7.13.0.564 (R2011b) NetCDF Library on 2013-05-08 14:45 UTC" ;
		:id = "ru29-20130507T211956" ;
		:institution = "Institute of Marine & Coastal Sciences, Rutgers University" ;
		:keywords = "Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "This data may be redistributed and used without restriction." ;
		:metadata_link = "" ;
		:naming_authority = "edu.rutgers.marine" ;
		:processing_level = "Dataset taken from glider native file format" ;
		:project = "Deployment not project based" ;
		:publisher_email = "kerfoot@marine.rutgers.edu" ;
		:publisher_name = "John Kerfoot" ;
		:publisher_url = "http://marine.rutgers.edu/cool/auvs" ;
		:sea_name = "" ;
		:standard_name_vocabulary = "CF-1.6" ;
		:summary = "The Rutgers University Coastal Ocean Observation Lab has deployed autonomous underwater gliders around the world since 1990.  Gliders are small, free-swimming, unmanned vehicles that use changes in buoyancy to move vertically and horizontally through the water column in a saw-tooth pattern.  They are deployed for days to several months and gather detailed information about the physical, chemical and biological processes of the world\'s  The Slocum glider was designed and oceans. built by Teledyne Webb Research Corporation, Falmouth, MA, USA." ;
		:time_coverage_end = "2013-05-08 07:56 UTC" ;
		:time_coverage_resolution = "point" ;
		:time_coverage_start = "2013-05-07 21:19 UTC" ;
		:title = "Slocum Glider Dataset" ;
}
