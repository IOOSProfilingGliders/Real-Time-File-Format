// Creator: kerfoot@marine.rutgers.edu
// Creation Date: 2013-05-09 15:00 EDT
// Common Data Language template for describing glider data using the
// Trajectory type.
//
// In addition to required global attributes, variables and variable
// attributes, this template does the following:
// 1. Creates a platform variable, where the name of the variable is one of:
//      slocum
//      seaglider
//      spray
//
//    This is an attempt to provide a means of identification of the glider
//    type which the NetCDF file originated from as there may be a need for
//    the DAC to do additional processing of the operator provided NetCDF 
//    files to bring them into compliance with the IOOS specification.
//
// 2. Addition of 2 new variables: segment_id and profile_id to identify the
//      underwater segment from the data was obtained.  As long as these are
//      sequentially numbered, it provides a means for the operators to
//      include multiple underwater segments, defined as the time between
//      surfacings, to include multiple segments in a single file.  Both
//      variables are dimensioned using the time coordinate variable and are
//      arrays containing an integer identifying the sequential segment
//      numbers.
//
// 3. Creation of 2 new variables: u and v.  These variables hold the
//      eastward_sea_water_velocity and northward_sea_water_velocity values
//      calculated by the glider during a segment, dive or profile.  They are
//      dimensioned using the trajectory coordinate as this made the most
//      sense since a single current is calculated for each segment, dive or
//      profile.  Not sure if this convention conforms to the CF Discrete 
//      Sampling Geometry guidelines or not.
//
// 4. Creation of 2 new qc variables: u_qc and v_qc.  Status flag variables
//      for specifying quality of the u and v values.
//
// 5. Addition of a global file attribute: netcdf_template_version.  Used to
//      track the evolution of the file specification.
//
// 7 General Variable Types:
//  COORDINATE
//  GEOSPATIAL
//  GEOPHYSICAL
//  ENUMERATED FLAG: geophysical variable qc flags
//  TRAJECTORY METADATA
//  PLATFORM
//  INSTRUMENT
netcdf glider_template {
dimensions:
	trajectory = 1 ;
	time = 1076 ;
variables:

    // COORDINATE variable enumerating the trajectory.
	int trajectory(trajectory) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:coordinates = "trajectory" ;
		trajectory:long_name = "Trajectory Name" ;

    // COORDINATE variable used to dimension all GEOSPATIAL, GEOPHYSICAL,
    // STATUS and TRAJECTORY METDATA variables
	double time(time) ;
		time:axis = "T" ;
		time:calendar = "gregorian" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;

    // TRAJECTORY METADATA variable
	int segment_id(time) ;
		segment_id:_FillValue = -2147483647 ;
        segment_id:comment = "Sequential segment number for the trajectory.  A segment is defined the collection of profiles contained in the trajectory" ;
		segment_id:long_name = "Segment ID" ;
		segment_id:valid_min = 1 ;
		segment_id:valid_max = 999 ;
		segment_id:observation_type = "calculated" ;
        segment_id:ancillary_variables = "platform profile_id trajectory" ;
        segment_id:platform = "platform" ;

    // TRAJECTORY METADATA variable
	int profile_id(time) ;
		profile_id:_FillValue = -2147483647 ;
        profile_id:comment = "Sequential profile number contained in the trajectory.  A profile is defined a single dive or climb" ;
		profile_id:long_name = "Profile ID" ;
		profile_id:valid_min = 1 ;
		profile_id:valid_max = 999 ;
		profile_id:observation_type = "calculated" ;
        profile_id:ancillary_variables = "platform segment_id trajectory" ;
        profile_id:platform = "platform" ;

    // GEOSPATIAL variable
	double depth(time) ;
		depth:_FillValue = 9.96920996838687e+36 ;
		depth:axis = "Z" ;
		depth:units = "meters" ;
		depth:standard_name = "depth" ;
		depth:valid_min = 0. ;
		depth:valid_max = 2000. ;
		depth:long_name = "Depth" ;
		depth:reference_datum = "sea-surface" ;
		depth:vertical_positive = "down" ;
		depth:observation_type = "calculated" ;
        depth:ancillary_variables = "depth_qc instrument_ctd" ;
        depth:platform = "platform" ;
        depth:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte depth_qc(time) ;
		depth_qc:_FillValue = -127b ;
		depth_qc:long_name = "depth Quality" ;
        depth:standard_name = "depth status_flag" ;
		depth_qc:flag_meanings =  ;
		depth_qc:valid_range = 0., 128. ;
		depth_qc:flag_values =  ;
        depth_qc:ancillary_variables = "depth instrument_ctd" ;

    // GEOSPATIAL variable
	double lat(time) ;
		lat:_FillValue = 9.96920996838687e+36 ;
		lat:axis = "Y" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
		lat:long_name = "Latitude" ;
		lat:observation_type = "measured" ;
        lat:ancillary_variables = "lat_qc" ;
        lat:platform = "platform" ;
    // ENUMERATED FLAG variable
	byte lat_qc(time) ;
		lat_qc:_FillValue = -127b ;
		lat_qc:long_name = "lat Quality" ;
        lat:standard_name = "lat status_flag" ;
		lat_qc:flag_meanings =  ;
		lat_qc:valid_range = 0., 128. ;
		lat_qc:flag_values =  ;
        lat_qc:ancillary_variables = "lat" ;

    // GEOSPATIAL variable
	double lon(time) ;
		lon:_FillValue = 9.96920996838687e+36 ;
		lon:axis = "X" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:long_name = "Longitude" ;
		lon:observation_type = "measured" ;
        lon:ancillary_variables = "lon" ;
        lon:platform = "platform" ;
    // ENUMERATED FLAG variable
	byte lon_qc(time) ;
		lon_qc:_FillValue = -127b ;
		lon_qc:long_name = "lon Quality" ;
        lon_qc:standard_name = "lon status_flag" ;
		lon_qc:flag_meanings =  ;
		lon_qc:valid_range = 0., 128. ;
		lon_qc:flag_values =  ;
        lon_qc:ancillary_variables = "lon" ;

    // GEOSPATIAL variable
	double pressure(time) ;
		pressure:_FillValue = 9.96920996838687e+36 ;
		pressure:axis = "Z" ;
		pressure:units = "dbar" ;
		pressure:standard_name = "pressure" ;
		pressure:valid_min = 0. ;
		pressure:valid_max = 2000. ;
		pressure:long_name = "Pressure" ;
		pressure:reference_datum = "sea-surface" ;
		pressure:vertical_positive = "down" ;
		pressure:observation_type = "measured" ;
        pressure:ancillary_variables = "pressure_qc instrument_ctd" ;
        pressure:platform = "platform" ;
        pressure:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte pressure_qc(time) ;
		pressure_qc:_FillValue = -127b ;
		pressure_qc:long_name = "pressure Quality" ;
        pressure_qc:standard_name = "pressure status_flag" ;
		pressure_qc:flag_meanings =  ;
		pressure_qc:valid_range = 0., 128. ;
		pressure_qc:flag_values =  ;
        pressure_qc:ancillary_variables = "pressure instrument_ctd" ;

    // GEOPHYSICAL variable
	double conductivity(time) ;
		conductivity:_FillValue = 9.96920996838687e+36 ;
		conductivity:units = "S m-1" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:valid_min = 0. ;
		conductivity:valid_max = 10. ;
		conductivity:long_name = "Sea Water Conductivity" ;
		conductivity:observation_type = "measured" ;
		conductivity:coordinates = "lon lat depth time" ;
        conductivity:ancillary_variables = "conductivity_qc instrument_ctd" ;
        conductivity:platform = "platform" ;
        conductivity:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte conductivity_qc(time) ;
		conductivity_qc:_FillValue = -127b ;
		conductivity_qc:long_name = "conductivity Quality" ;
        conductivity_qc:standard_name = "conductivity status_flag" ;
		conductivity_qc:flag_meanings =  ;
		conductivity_qc:valid_range = 0., 128. ;
		conductivity_qc:flag_values =  ;
        conductivity:ancillary_variables = "conductivity instrument_ctd" ;

    // GEOPHYSICAL variable
	double density(time) ;
		density:_FillValue = 9.96920996838687e+36 ;
		density:units = "kg m-3" ;
		density:standard_name = "sea_water_density" ;
		density:valid_min = 1015. ;
		density:valid_max = 1040. ;
		density:long_name = "Sea Water Density" ;
		density:observation_type = "calculated" ;
		density:coordinates = "lon lat depth time" ;
        density:ancillary_variables = "density_qc instrument_ctd" ;
        density:platform = "platform" ;
        density:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte density_qc(time) ;
		density_qc:_FillValue = -127b ;
		density_qc:long_name = "density Quality" ;
        density_qc:standard_name = "density status_flag" ;
		density_qc:flag_meanings =  ;
		density_qc:valid_range = 0., 128. ;
		density_qc:flag_values =  ;
        density_qc:ancillary_variables = "density instrument_ctd" ;

    // GEOPHYSICAL variable
	double salinity(time) ;
		salinity:_FillValue = 9.96920996838687e+36 ;
		salinity:units = "1e-3" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:valid_min = 0. ;
		salinity:valid_max = 40. ;
		salinity:long_name = "Sea Water Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:coordinates = "lon lat depth time" ;
        salinity:ancillary_variables = "salinity_qc instrument_ctd" ;
        salinity:platform = "platform" ;
        salinity:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte salinity_qc(time) ;
		salinity_qc:_FillValue = -127b ;
		salinity_qc:long_name = "salinity Quality" ;
        salinity_qc:standard_name = "salinity status_flag" ;
		salinity_qc:flag_meanings =  ;
		salinity_qc:valid_range = 0., 128. ;
		salinity_qc:flag_values =  ;
        salinity_qc:ancillary_variables = "salinity instrument_ctd" ;

    // GEOPHYSICAL variable
	double temperature(time) ;
		temperature:_FillValue = 9.96920996838687e+36 ;
		temperature:units = "Celsius" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:valid_min = -5. ;
		temperature:valid_max = 40. ;
		temperature:long_name = "Sea Water Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:coordinates = "lon lat depth time" ;
        temperature:ancillary_variables = "temperature_qc instrument_ctd" ;
        temperature:platform = "platform" ;
        temperature:instrument = "instrument_ctd" ;
    // ENUMERATED FLAG variable
	byte temperature_qc(time) ;
		temperature_qc:_FillValue = -127b ;
		temperature_qc:long_name = "temperature Quality" ;
        temperature_qc:standard_name = "temperature status_flag" ;
		temperature_qc:flag_meanings =  ;
		temperature_qc:valid_range = 0., 128. ;
		temperature_qc:flag_values =  ;
        temperature_qc:ancillary_variables = "temperature instrument_ctd" ;

	double u(trajectory) ;
		u:_FillValue = 9.96920996838687e+36 ;
		u:units = "m s-1" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:valid_min = 0. ;
		u:valid_max = 3. ;
		u:long_name = "Eastward Sea Water Velocity" ;
		u:observation_type = "calculated" ;
		u:coordinates = "trajectory" ;
	byte u_qc(trajectory) ;
		u_qc:_FillValue = -127b ;
		u_qc:long_name = "u Quality" ;
		u_qc:flag_meanings =  ;
		u_qc:valid_range = 0., 128. ;
		u_qc:flag_values =  ;

	double v(trajectory) ;
		v:_FillValue = 9.96920996838687e+36 ;
		v:units = "m s-1" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:valid_min = 0. ;
		v:valid_max = 3. ;
		v:long_name = "Northward Sea Water Velocity" ;
		v:observation_type = "calculated" ;
		v:coordinates = "trajectory" ;

	byte v_qc(trajectory) ;
		v_qc:_FillValue = -127b ;
		v_qc:long_name = "v Quality" ;
		v_qc:flag_meanings =  ;
		v_qc:valid_range = 0., 128. ;
		v_qc:flag_values =  ;

    // PLATFORM variable
	int slocum ;
		platform:wmo_id = "ru29" ;
		platform:comment = "Slocum Glider ru29" ;
		platform:id = "ru29" ;
		platform:long_name = "Slocum Glider ru29" ;

    // INSTRUMENT variable
	int instrument_ctd ;
		instrument_ctd:comment = "Unpumped CTD with a nominal sampling rate of 1Hz." ;
		instrument_ctd:serial_number =  ;
		instrument_ctd:long_name = "Seabird SBD 41CP Conductivity, Temperature, Depth Sensor." ;
        instrument_ctd:ancillary_variables = "platform temperature temperature_qc salinity salinity_qc pressure pressure_qc depth depth_qc conductivity conductivity_qc"

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:acknowledgment =  ;
		:cdm_data_type = "Trajectory" ;
		:comment =  ;
		:contributor_name = "Scott Glenn, Oscar Schofield, John Kerfoot" ;
		:contributor_role = "Principal Investigator, Principal Investigator, Data Manager" ;
		:creator_email = "kerfoot@marine.rutgers.edu" ;
		:creator_name = "John Kerfoot" ;
		:creator_url = "http://marine.rutgers.edu/cool/auvs" ;
		:date_created = "2013-05-08 14:45 UTC" ;
		:date_issued = "2013-05-08 14:45 UTC" ;
		:date_modified = "2013-05-08 14:45 UTC" ;
		:featureType = "trajectory" ;
        // file_version attribute to track changes in the template
        :netcdf_template_version = "IOOS_Glider_NetCDF_Trajectory_Template_v1.0" ;
		:geospatial_lat_max = -15.88833 ;
		:geospatial_lat_min = -15.9445416666667 ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 1.49547333333333 ;
		:geospatial_lon_min = 1.394655 ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_max = 987.26 ;
		:geospatial_vertical_min = 0. ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_units = "meters" ;
		:history = "Created with the Matlab 7.13.0.564 (R2011b) NetCDF Library on 2013-05-08 14:45 UTC" ;
		:id = "ru29-20130507T211956" ;
		:institution = "Institute of Marine & Coastal Sciences, Rutgers University" ;
		:keywords = "Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "This data may be redistributed and used without restriction." ;
		:metadata_link =  ;
		:naming_authority = "edu.rutgers.marine" ;
		:processing_level = "Dataset taken from glider native file format" ;
		:project = "Deployment not project based" ;
		:publisher_email = "kerfoot@marine.rutgers.edu" ;
		:publisher_name = "John Kerfoot" ;
		:publisher_url = "http://marine.rutgers.edu/cool/auvs" ;
		:sea_name =  ;
		:standard_name_vocabulary = "CF-1.6" ;
		:summary = "The Rutgers University Coastal Ocean Observation Lab has deployed autonomous underwater gliders around the world since 1990.  Gliders are small, free-swimming, unmanned vehicles that use changes in buoyancy to move vertically and horizontally through the water column in a saw-tooth pattern.  They are deployed for days to several months and gather detailed information about the physical, chemical and biological processes of the world\'s  The Slocum glider was designed and oceans. built by Teledyne Webb Research Corporation, Falmouth, MA, USA." ;
		:time_coverage_end = "2013-05-08 07:56 UTC" ;
		:time_coverage_resolution = "point" ;
		:time_coverage_start = "2013-05-07 21:19 UTC" ;
		:title = "Slocum Glider Dataset" ;
}
