netcdf glider_trajectory_uv_template_v.0.0 {
dimensions:
	time = UNLIMITED ; // (0 currently)
	trajectory = 1 ;
	time_uv = 1 ;
variables:
	double time(time) ;
		time:axis = "T" ;
		time:calendar = "gregorian" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;
		time:sensor_name =  ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
	byte time_qc(time) ;
		time_qc:_FillValue = -127b ;
		time_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		time_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		time_qc:long_name = "time Quality Flag" ;
		time_qc:standard_name = "time status_flag" ;
		time_qc:valid_max = 9b ;
		time_qc:valid_min = 0b ;
	double time_uv(time_uv) ;
		time_uv:axis = "T" ;
		time_uv:calendar = "gregorian" ;
		time_uv:long_name = "Approximate time midpoint of each segment" ;
		time_uv:observation_type = "estimated" ;
		time_uv:standard_name = "time" ;
		time_uv:units = "seconds since 1970-01-01 00:00:00 UTC" ;
	short trajectory(trajectory) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "A trajectory can span multiple data files each containing a single segment." ;
		trajectory:long_name = "Unique identifier for each trajectory feature contained in the file" ;
	short segment_id(time) ;
		segment_id:_FillValue = -32767s ;
		segment_id:comment = "Sequential segment number within a trajectory/deployment. A segment corresponds to the set of data collected between 2 gps fixes obtained when the glider surfaces." ;
		segment_id:long_name = "Segment ID" ;
		segment_id:observation_type = "calculated" ;
		segment_id:valid_max = 999 ;
		segment_id:valid_min = 1 ;
	short profile_id(time) ;
		profile_id:_FillValue = -32767s ;
		profile_id:comment = "Sequential profile number within the current segment. A profile is defined as a single dive or climb" ;
		profile_id:long_name = "Profile ID" ;
		profile_id:observation_type = "calculated" ;
		profile_id:valid_max = 999 ;
		profile_id:valid_min = 1 ;
	double depth(time) ;
		depth:_FillValue = 9.96920996838687e+36 ;
		depth:ancillary_variables = "depth_qc" ;
		depth:axis = "Z" ;
		depth:instrument = "instrument_ctd" ;
		depth:long_name = "Depth" ;
		depth:observation_type = "calculated" ;
		depth:platform = "platform" ;
		depth:positive = "down" ;
		depth:reference_datum = "sea-surface" ;
		depth:sensor_name =  ;
		depth:standard_name = "depth" ;
		depth:units = "meters" ;
		depth:valid_max = 2000 ;
		depth:valid_min = 0 ;
	byte depth_qc(time) ;
		depth_qc:_FillValue = -127b ;
		depth_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		depth_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		depth_qc:long_name = "depth Quality Flag" ;
		depth_qc:standard_name = "depth status_flag" ;
		depth_qc:valid_max = 9b ;
		depth_qc:valid_min = 0b ;
	double lat(time) ;
		lat:_FillValue = 9.96920996838687e+36 ;
		lat:ancillary_variables = "lat_qc" ;
		lat:axis = "Y" ;
		lat:comment = "Some values are linearly interpolated between measured coordinates.  See lat_qc" ;
		lat:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lat:flag_meanings =  ;
		lat:long_name = "Latitude" ;
		lat:observation_type = "measured" ;
		lat:platform = "platform" ;
		lat:reference = "WGS84" ;
		lat:sensor_name =  ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
	byte lat_qc(time) ;
		lat_qc:_FillValue = -127b ;
		lat_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		lat_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lat_qc:long_name = "lat Quality Flag" ;
		lat_qc:standard_name = "lat status_flag" ;
		lat_qc:valid_max = 9b ;
		lat_qc:valid_min = 0b ;
	double lon(time) ;
		lon:_FillValue = 9.96920996838687e+36 ;
		lon:ancillary_variables = "lon_qc" ;
		lon:axis = "X" ;
		lon:comment = "Some values are linearly interpolated between measured coordinates.  See lon_qc" ;
		lon:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lon:flag_meanings =  ;
		lon:long_name = "Longitude" ;
		lon:observation_type = "measured" ;
		lon:platform = "platform" ;
		lon:reference = "WGS84" ;
		lon:sensor_name =  ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
	byte lon_qc(time) ;
		lon_qc:_FillValue = -127b ;
		lon_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		lon_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lon_qc:long_name = "lon Quality Flag" ;
		lon_qc:standard_name = "lon status_flag" ;
		lon_qc:valid_max = 9b ;
		lon_qc:valid_min = 0b ;
	double pressure(time) ;
		pressure:_FillValue = 9.96920996838687e+36 ;
		pressure:accuracy =  ;
		pressure:ancillary_variables = "pressure_qc" ;
		pressure:axis = "Z" ;
		pressure:instrument = "instrument_ctd" ;
		pressure:long_name = "Pressure" ;
		pressure:observation_type = "calculated" ;
		pressure:platform = "platform" ;
		pressure:positive = "down" ;
		pressure:precision =  ;
		pressure:reference_datum = "sea-surface" ;
		pressure:resolution =  ;
		pressure:sensor_name =  ;
		pressure:standard_name = "pressure" ;
		pressure:units = "dbar" ;
		pressure:valid_max = 2000 ;
		pressure:valid_min = 0 ;
	byte pressure_qc(time) ;
		pressure_qc:_FillValue = -127b ;
		pressure_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		pressure_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		pressure_qc:long_name = "pressure Quality Flag" ;
		pressure_qc:standard_name = "pressure status_flag" ;
		pressure_qc:valid_max = 9b ;
		pressure_qc:valid_min = 0b ;
	double conductivity(time) ;
		conductivity:_FillValue = 9.96920996838687e+36 ;
		conductivity:accuracy =  ;
		conductivity:ancillary_variables = "conductivity_qc" ;
		conductivity:coordinates = "lon lat depth time" ;
		conductivity:instrument = "instrument_ctd" ;
		conductivity:long_name = "Conductivity" ;
		conductivity:observation_type = "measured" ;
		conductivity:platform = "platform" ;
		conductivity:precision =  ;
		conductivity:resolution =  ;
		conductivity:sensor_name =  ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:valid_max = 10. ;
		conductivity:valid_min = 0. ;
	byte conductivity_qc(time) ;
		conductivity_qc:_FillValue = -127b ;
		conductivity_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		conductivity_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		conductivity_qc:long_name = "conductivity Quality Flag" ;
		conductivity_qc:standard_name = "conductivity status_flag" ;
		conductivity_qc:valid_max = 9b ;
		conductivity_qc:valid_min = 0b ;
	double density(time) ;
		density:_FillValue = 9.96920996838687e+36 ;
		density:ancillary_variables = "density_qc" ;
		density:coordinates = "lon lat depth time" ;
		density:instrument = "instrument_ctd" ;
		density:long_name = "Density" ;
		density:observation_type = "calculated" ;
		density:platform = "platform" ;
		density:sensor_name =  ;
		density:standard_name = "sea_water_density" ;
		density:units = "kg m-3" ;
		density:valid_max = 1040. ;
		density:valid_min = 1015. ;
	byte density_qc(time) ;
		density_qc:_FillValue = -127b ;
		density_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		density_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		density_qc:long_name = "density Quality Flag" ;
		density_qc:standard_name = "density status_flag" ;
		density_qc:valid_max = 9b ;
		density_qc:valid_min = 0b ;
	double salinity(time) ;
		salinity:_FillValue = 9.96920996838687e+36 ;
		salinity:ancillary_variables = "salinity_qc" ;
		salinity:coordinates = "lon lat depth time" ;
		salinity:instrument = "instrument_ctd" ;
		salinity:long_name = "Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:platform = "platform" ;
		salinity:sensor_name =  ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:units = "1e-3" ;
		salinity:valid_max = 40. ;
		salinity:valid_min = 0. ;
	byte salinity_qc(time) ;
		salinity_qc:_FillValue = -127b ;
		salinity_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		salinity_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		salinity_qc:long_name = "salinity Quality Flag" ;
		salinity_qc:standard_name = "salinity status_flag" ;
		salinity_qc:valid_max = 9b ;
		salinity_qc:valid_min = 0b ;
	double temperature(time) ;
		temperature:_FillValue = 9.96920996838687e+36 ;
		temperature:accuracy =  ;
		temperature:ancillary_variables = "temperature_qc" ;
		temperature:coordinates = "lon lat depth time" ;
		temperature:instrument = "instrument_ctd" ;
		temperature:long_name = "Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:platform = "platform" ;
		temperature:precision =  ;
		temperature:resolution =  ;
		temperature:sensor_name =  ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:valid_max = 40. ;
		temperature:valid_min = -5. ;
	byte temperature_qc(time) ;
		temperature_qc:_FillValue = -127b ;
		temperature_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		temperature_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		temperature_qc:long_name = "temperature Quality Flag" ;
		temperature_qc:standard_name = "temperature status_flag" ;
		temperature_qc:valid_max = 9b ;
		temperature_qc:valid_min = 0b ;
	double lat_uv(time_uv) ;
		lat_uv:_FillValue = 9.96920996838687e+36 ;
		lat_uv:axis = "Y" ;
		lat_uv:comment = "Values are interpolated to provide the center latitude of the segment" ;
		lat_uv:long_name = "Center Latitude for Depth-Averaged Current" ;
		lat_uv:observation_type = "calculated" ;
		lat_uv:platform = "platform" ;
		lat_uv:standard_name = "latitude" ;
		lat_uv:units = "degrees_north" ;
		lat_uv:valid_max = 90. ;
		lat_uv:valid_min = -90. ;
	double lon_uv(time_uv) ;
		lon_uv:_FillValue = 9.96920996838687e+36 ;
		lon_uv:axis = "X" ;
		lon_uv:comment = "Values are interpolated to provide the center longitude of the segment" ;
		lon_uv:long_name = "Center Longitude for Depth-Averaged Current" ;
		lon_uv:observation_type = "calculated" ;
		lon_uv:platform = "platform" ;
		lon_uv:standard_name = "longitude" ;
		lon_uv:units = "degrees_east" ;
		lon_uv:valid_max = 180. ;
		lon_uv:valid_min = -180. ;
	double u(time_uv) ;
		u:_FillValue = 9.96920996838687e+36 ;
		u:coordinates = "lon_uv lat_uv time_uv" ;
		u:long_name = "Eastward Sea Water Velocity" ;
		u:observation_type = "calculated" ;
		u:platform = "platform" ;
		u:sensor_name =  ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:units = "m s-1" ;
		u:valid_max = 10. ;
		u:valid_min = -10. ;
	byte u_qc(time_uv) ;
		u_qc:_FillValue = -127b ;
		u_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		u_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		u_qc:long_name = "u Quality Flag" ;
		u_qc:standard_name = "u status_flag" ;
		u_qc:valid_max = 9b ;
		u_qc:valid_min = 0b ;
	double v(time_uv) ;
		v:_FillValue = 9.96920996838687e+36 ;
		v:coordinates = "lon_uv lat_uv time_uv" ;
		v:long_name = "Northward Sea Water Velocity" ;
		v:observation_type = "calculated" ;
		v:platform = "platform" ;
		v:sensor_name =  ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:units = "m s-1" ;
		v:valid_max = 10. ;
		v:valid_min = -10. ;
	byte v_qc(time_uv) ;
		v_qc:_FillValue = -127b ;
		v_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed interpolated_value missing_value" ;
		v_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		v_qc:long_name = "v Quality Flag" ;
		v_qc:standard_name = "v status_flag" ;
		v_qc:valid_max = 9b ;
		v_qc:valid_min = 0b ;
	byte platform ;
		platform:comment = "Slocum Glider ru29" ;
		platform:id = "ru29" ;
		platform:instrument = "instrument_ctd" ;
		platform:long_name = "Slocum Glider ru29" ;
		platform:type = "platform" ;
		platform:wmo_id = "ru29" ;
	byte instrument_ctd ;
		instrument_ctd:calibration_date = "2000-01-01" ;
		instrument_ctd:calibration_report =  ;
		instrument_ctd:comment = "Slocum Glider ru29" ;
		instrument_ctd:factory_calibrated =  ;
		instrument_ctd:long_name = "Seabird SBD 41CP Conductivity, Temperature, Depth Sensor" ;
		instrument_ctd:make_model = "Seabird SBE 41CP" ;
		instrument_ctd:platform = "platform" ;
		instrument_ctd:serial_number = "0098" ;
		instrument_ctd:user_calibrated =  ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:acknowledgment = "This deployment partially supported by ..." ;
		:cdm_data_type = "Trajectory" ;
		:comment = "This file is intended to be used as a template only.  Data is not to be used for scientific purposes." ;
		:contributor_name = "Scott Glenn, Oscar Schofield, John Kerfoot" ;
		:contributor_role = "Principal Investigator, Principal Investigator, Data Manager" ;
		:creator_email = "kerfoot@marine.rutgers.edu" ;
		:creator_name = "John Kerfoot" ;
		:creator_url = "http://marine.rutgers.edu/cool/auvs" ;
		:date_created = "2013-05-08 14:45 UTC" ;
		:date_issued = "2013-05-08 14:45 UTC" ;
		:date_modified = "2013-05-08 14:45 UTC" ;
		:featureType = "trajectory" ;
		:format_version = "IOOS_Glider_NetCDF_Trajectory_Template_v0.0" ;
		:geospatial_lat_max = -15.88833 ;
		:geospatial_lat_min = -15.9445416666667 ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_max = 1.49547333333333 ;
		:geospatial_lon_min = 1.394655 ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_max = 987.26 ;
		:geospatial_vertical_min = 0. ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_units = "meters" ;
		:history = "Created on Wed Aug  7 07:27:21 2013" ;
		:id = "ru29-20130507T211956" ;
		:institution = "Institute of Marine & Coastal Sciences, Rutgers University" ;
		:keywords = "Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "This data may be redistributed and used without restriction." ;
		:metadata_link =  ;
		:naming_authority = "edu.rutgers.marine" ;
		:processing_level = "Dataset taken from glider native file format" ;
		:project = "Deployment not project based" ;
		:publisher_email = "kerfoot@marine.rutgers.edu" ;
		:publisher_name = "John Kerfoot" ;
		:publisher_url = "http://marine.rutgers.edu/cool/auvs" ;
		:references =  ;
		:sea_name = "South Atlantic Ocean" ;
		:source = "Observational data from a profiling glider" ;
		:standard_name_vocabulary = "CF-v25" ;
		:summary = "The Rutgers University Coastal Ocean Observation Lab has deployed autonomous underwater gliders around the world since 1990. Gliders are small, free-swimming, unmanned vehicles that use changes in buoyancy to move vertically and horizontally through the water column in a saw-tooth pattern. They are deployed for days to several months and gather detailed information about the physical, chemical and biological processes of the world\'s The Slocum glider was designed and oceans. built by Teledyne Webb Research Corporation, Falmouth, MA, USA." ;
		:time_coverage_end = "2013-05-08 07:56 UTC" ;
		:time_coverage_resolution = "point" ;
		:time_coverage_start = "2013-05-07 21:19 UTC" ;
		:title = "Slocum Glider Dataset" ;
}
