netcdf C:/Users/derrick.snowden/Documents/GitHub/Real-Time-File-Format/examples/proposed_templates/glider_trajectory_uv_template_v.0.0.nc {
 dimensions:
   time = UNLIMITED;   // (0 currently)
   time_uv = 1;
   trajectory = 1;
 variables:
   double time(time=0);
     :axis = "T";
     :calendar = "gregorian";
     :long_name = "Time";
     :observation_type = "measured";
     :standard_name = "time";
     :units = "seconds since 1970-01-01 00:00:00 UTC";
     :_ChunkSize = 1; // int
   double time_uv(time_uv=1);
     :axis = "T";
     :calendar = "gregorian";
     :long_name = "Approximate time midpoint of each segment";
     :observation_type = "estimated";
     :standard_name = "time";
     :units = "seconds since 1970-01-01 00:00:00 UTC";
     :_ChunkSize = 1; // int
   short trajectory(trajectory=1);
     :cf_role = "trajectory_id";
     :comment = "A trajectory can span multiple data files each containing a single segment.";
     :long_name = "Unique identifier for each trajectory feature contained in the file";
     :_ChunkSize = 1; // int
   short segment_id(time=0);
     :comment = "Sequential segment number within a trajectory/deployment. A segment corresponds to the set of data collected between 2 gps fixes obtained when the glider surfaces.";
     :long_name = "Segment ID";
     :observation_type = "calculated";
     :valid_max = 999; // int
     :valid_min = 1; // int
     :_FillValue = -32767S; // short
     :_ChunkSize = 1; // int
   short profile_id(time=0);
     :_FillValue = -32767S; // short
     :comment = "Sequential profile number within the current segment. A profile is defined as a single dive or climb";
     :long_name = "Profile ID";
     :observation_type = "calculated";
     :valid_max = 999; // int
     :valid_min = 1; // int
     :_ChunkSize = 1; // int
   double depth(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "depth_qc";
     :axis = "Z";
     :instrument = "instrument_ctd";
     :long_name = "Depth";
     :observation_type = "calculated";
     :platform = "platform";
     :positive = "down";
     :reference_datum = "sea-surface";
     :standard_name = "depth";
     :units = "meters";
     :valid_max = 2000; // int
     :valid_min = 0; // int
     :_ChunkSize = 1; // int
   byte depth_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "depth Quality Flag";
     :standard_name = "depth status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double lat(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "lat_qc";
     :axis = "Y";
     :comment = "Some values are linearly interpolated between measured coordinates.  See lat_qc";
     :flag_meanings = "";
     :long_name = "Latitude";
     :observation_type = "measured";
     :platform = "platform";
     :standard_name = "latitude";
     :units = "degrees_north";
     :valid_max = 90.0; // double
     :valid_min = -90.0; // double
     :_ChunkSize = 1; // int
   byte lat_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "lat Quality Flag";
     :standard_name = "lat status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double lon(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "lon_qc";
     :axis = "X";
     :comment = "Some values are linearly interpolated between measured coordinates.  See lon_qc";
     :flag_meanings = "";
     :long_name = "Longitude";
     :observation_type = "measured";
     :platform = "platform";
     :standard_name = "longitude";
     :units = "degrees_east";
     :valid_max = 180.0; // double
     :valid_min = -180.0; // double
     :_ChunkSize = 1; // int
   byte lon_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "lon Quality Flag";
     :standard_name = "lon status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double pressure(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "pressure_qc";
     :axis = "Z";
     :instrument = "instrument_ctd";
     :long_name = "Pressure";
     :observation_type = "calculated";
     :platform = "platform";
     :positive = "down";
     :reference_datum = "sea-surface";
     :standard_name = "pressure";
     :units = "dbar";
     :valid_max = 2000; // int
     :valid_min = 0; // int
     :_ChunkSize = 1; // int
   byte pressure_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "pressure Quality Flag";
     :standard_name = "pressure status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double conductivity(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "conductivity_qc";
     :coordinates = "lon lat depth time";
     :instrument = "instrument_ctd";
     :long_name = "Conductivity";
     :observation_type = "measured";
     :platform = "platform";
     :standard_name = "sea_water_electrical_conductivity";
     :units = "S m-1";
     :valid_max = 10.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   byte conductivity_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "conductivity Quality Flag";
     :standard_name = "conductivity status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double density(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "density_qc";
     :coordinates = "lon lat depth time";
     :instrument = "instrument_ctd";
     :long_name = "Density";
     :observation_type = "calculated";
     :platform = "platform";
     :standard_name = "sea_water_density";
     :units = "kg m-3";
     :valid_max = 1040.0; // double
     :valid_min = 1015.0; // double
     :_ChunkSize = 1; // int
   byte density_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "density Quality Flag";
     :standard_name = "density status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double salinity(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "salinity_qc";
     :coordinates = "lon lat depth time";
     :instrument = "instrument_ctd";
     :long_name = "Salinity";
     :observation_type = "calculated";
     :platform = "platform";
     :standard_name = "sea_water_salinity";
     :units = "1e-3";
     :valid_max = 40.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   byte salinity_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "salinity Quality Flag";
     :standard_name = "salinity status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double temperature(time=0);
     :_FillValue = 9.969209968386869E36; // double
     :ancillary_variables = "temperature_qc";
     :coordinates = "lon lat depth time";
     :instrument = "instrument_ctd";
     :long_name = "Temperature";
     :observation_type = "measured";
     :platform = "platform";
     :standard_name = "sea_water_temperature";
     :units = "Celsius";
     :valid_max = 40.0; // double
     :valid_min = -5.0; // double
     :_ChunkSize = 1; // int
   byte temperature_qc(time=0);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "temperature Quality Flag";
     :standard_name = "temperature status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double u(time_uv=1);
     :_FillValue = 9.969209968386869E36; // double
     :coordinates = "time_uv";
     :long_name = "Eastward Sea Water Velocity";
     :observation_type = "calculated";
     :platform = "platform";
     :standard_name = "eastward_sea_water_velocity";
     :units = "m s-1";
     :valid_max = 10.0; // double
     :valid_min = -10.0; // double
     :_ChunkSize = 1; // int
   byte u_qc(time_uv=1);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "u Quality Flag";
     :standard_name = "u status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   double v(time_uv=1);
     :_FillValue = 9.969209968386869E36; // double
     :coordinates = "time_uv";
     :long_name = "Northward Sea Water Velocity";
     :observation_type = "calculated";
     :platform = "platform";
     :standard_name = "northward_sea_water_velocity";
     :units = "m s-1";
     :valid_max = 10.0; // double
     :valid_min = -10.0; // double
     :_ChunkSize = 1; // int
   byte v_qc(time_uv=1);
     :_FillValue = -127B; // byte
     :flag_meanings = "";
     :flag_values = "";
     :long_name = "v Quality Flag";
     :standard_name = "v status_flag";
     :valid_max = 128.0; // double
     :valid_min = 0.0; // double
     :_ChunkSize = 1; // int
   byte platform;
     :comment = "Slocum Glider ru29";
     :id = "ru29";
     :instrument = "instrument_ctd";
     :long_name = "Slocum Glider ru29";
     :type = "platform";
     :wmo_id = "ru29";
   byte instrument_ctd;
     :accuracy = "";
     :calibration_date = "2000-01-01";
     :calibration_report = "";
     :comment = "Slocum Glider ru29";
     :factory_calibrated = "";
     :long_name = "Seabird SBD 41CP Conductivity, Temperature, Depth Sensor";
     :make_model = "Seabird SBE 41CP";
     :platform = "platform";
     :precision = "";
     :serial_number = "0098";
     :user_calibrated = "";
     :valid_range = "";

 :Conventions = "CF-1.6";
 :Metadata_Conventions = "Unidata Dataset Discovery v1.0";
 :acknowledgment = "This deployment partially supported by ...";
 :cdm_data_type = "Trajectory";
 :comment = "This file is intended to be used as a template only.  Data is not to be used for scientific purposes.";
 :contributor_name = "Scott Glenn, Oscar Schofield, John Kerfoot";
 :contributor_role = "Principal Investigator, Principal Investigator, Data Manager";
 :creator_email = "kerfoot@marine.rutgers.edu";
 :creator_name = "John Kerfoot";
 :creator_url = "http://marine.rutgers.edu/cool/auvs";
 :date_created = "2013-05-08 14:45 UTC";
 :date_issued = "2013-05-08 14:45 UTC";
 :date_modified = "2013-05-08 14:45 UTC";
 :featureType = "trajectory";
 :file_version = "IOOS_Glider_NetCDF_Trajectory_Template_v0.0";
 :geospatial_lat_max = -15.88833; // double
 :geospatial_lat_min = -15.9445416666667; // double
 :geospatial_lat_resolution = "point";
 :geospatial_lat_units = "degrees_north";
 :geospatial_lon_max = 1.49547333333333; // double
 :geospatial_lon_min = 1.394655; // double
 :geospatial_lon_resolution = "point";
 :geospatial_lon_units = "degrees_east";
 :geospatial_vertical_max = 987.26; // double
 :geospatial_vertical_min = 0.0; // double
 :geospatial_vertical_positive = "down";
 :geospatial_vertical_resolution = "point";
 :geospatial_vertical_units = "meters";
 :history = "Created on Mon Jul 22 15:49:44 2013";
 :id = "ru29-20130507T211956";
 :institution = "Institute of Marine & Coastal Sciences, Rutgers University";
 :keywords = "Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity";
 :keywords_vocabulary = "GCMD Science Keywords";
 :license = "This data may be redistributed and used without restriction.";
 :metadata_link = "";
 :naming_authority = "edu.rutgers.marine";
 :processing_level = "Dataset taken from glider native file format";
 :project = "Deployment not project based";
 :publisher_email = "kerfoot@marine.rutgers.edu";
 :publisher_name = "John Kerfoot";
 :publisher_url = "http://marine.rutgers.edu/cool/auvs";
 :references = "";
 :sea_name = "South Atlantic Ocean";
 :source = "Observational data from a profiling glider";
 :standard_name_vocabulary = "CF-v25";
 :summary = "The Rutgers University Coastal Ocean Observation Lab has deployed autonomous underwater gliders around the world since 1990. Gliders are small, free-swimming, unmanned vehicles that use changes in buoyancy to move vertically and horizontally through the water column in a saw-tooth pattern. They are deployed for days to several months and gather detailed information about the physical, chemical and biological processes of the world\'s The Slocum glider was designed and oceans. built by Teledyne Webb Research Corporation, Falmouth, MA, USA.";
 :time_coverage_end = "2013-05-08 07:56 UTC";
 :time_coverage_resolution = "point";
 :time_coverage_start = "2013-05-07 21:19 UTC";
 :title = "Slocum Glider Dataset";
}
